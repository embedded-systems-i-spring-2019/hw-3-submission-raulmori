fdfdfadf
